module layer1
