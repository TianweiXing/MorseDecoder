module rom();
  reg [31:0] inputs[0:25];
  reg [34:0] weights[0:30];
  initial begin
    inputs[0] =  32'b_00000000_00000000_00000011_00001001;
    inputs[1] =  32'b_00001001_00000011_00000011_00000011;
    inputs[2] =  32'b_00001001_00000011_00001001_00000011;
    inputs[3] =  32'b_00000000_00001001_00000011_00000011;
    inputs[4] =  32'b_00000000_00000000_00000000_00000011;
    inputs[5] =  32'b_00000011_00000011_00001001_00000011;
    inputs[6] =  32'b_00000000_00001001_00001001_00000011;
    inputs[7] =  32'b_00000011_00000011_00000011_00000011;
    inputs[8] =  32'b_00000000_00000000_00000011_00000011;
    inputs[9] =  32'b_00000011_00001001_00001001_00001001;
    inputs[10] =  32'b_00000000_00001001_00000011_00001001;
    inputs[11] =  32'b_00000011_00001001_00000011_00000011;
    inputs[12] =  32'b_00000000_00000000_00001001_00001001;
    inputs[13] =  32'b_00000000_00000000_00001001_00000011;
    inputs[14] =  32'b_00000000_00001001_00001001_00001001;
    inputs[15] =  32'b_00000011_00001001_00001001_00000011;
    inputs[16] =  32'b_00001001_00001001_00000011_00001001;
    inputs[17] =  32'b_00000000_00000011_00001001_00000011;
    inputs[18] =  32'b_00000000_00000011_00000011_00000011;
    inputs[19] =  32'b_00000000_00000000_00000000_00001001;
    inputs[20] =  32'b_00000000_00000011_00000011_00001001;
    inputs[21] =  32'b_00000011_00000011_00000011_00001001;
    inputs[22] =  32'b_00000000_00000011_00001001_00001001;
    inputs[23] =  32'b_00001001_00000011_00000011_00001001;
    inputs[24] =  32'b_00001001_00000011_00001001_00001001;
    inputs[25] =  32'b_00001001_00001001_00000011_00000011;

    weights[0] =  35'b_0010011_0001001_1111110_0000101_1111000;
    weights[1] =  35'b_1111010_0000001_1111101_1111100_0000001;
    weights[2] =  35'b_0001010_1101100_0001001_0010000_0001000;
    weights[3] =  35'b_0001010_1110101_0011110_0001111_1011101;

    weights[4] =  35'b_1110000_0000001_0010011_1111101_1101100;
    weights[5] =  35'b_0001011_0000011_0001100_1110011_0000110;
    weights[6] =  35'b_0000000_1111111_1111011_0000111_1101001;
    weights[7] =  35'b_0010000_0000000_1110110_1011100_0010010;
    weights[8] =  35'b_1110001_1111101_0011011_1101111_0010111;
    weights[9] =  35'b_1111000_0000101_1111001_0001100_1100110;
    weights[10] =  35'b_1110111_0000001_1100000_0010001_0001110;
    weights[11] =  35'b_0000101_0000010_0000000_0000000_0011100;
    weights[12] =  35'b_1100000_1111101_0010000_0000000_0011100;
    weights[13] =  35'b_0000101_1111110_1110000_0001001_1100110;
    weights[14] =  35'b_0000110_0000000_1101000_0000111_0100001;
    weights[15] =  35'b_0001101_0000100_0000000_1110101_0001000;
    weights[16] =  35'b_1101101_0000010_0001010_0000100_1101100;
    weights[17] =  35'b_1100111_0000010_0000000_0001010_0001001;
    weights[18] =  35'b_1111001_1111101_1101011_0010000_1101110;
    weights[19] =  35'b_0000011_1111111_1100111_0001100_1101111;
    weights[20] =  35'b_0001011_1111101_1111110_1111101_1101000;
    weights[21] =  35'b_1110010_0000001_1110000_0010000_1110110;
    weights[22] =  35'b_1111110_0000000_1110101_0001010_0101000;
    weights[23] =  35'b_1111010_0000011_0010111_1110111_1110010;
    weights[24] =  35'b_1110110_0000011_0001010_0000010_0010100;
    weights[25] =  35'b_0000001_1111010_0001101_1111011_0000001;
    weights[26] =  35'b_1110100_0000111_0000010_0001000_1110010;
    weights[27] =  35'b_0000111_0000100_0010101_1110001_1100110;
    weights[28] =  35'b_1111101_1111011_0000101_0000011_1101101;
    weights[29] =  35'b_0001010_0000011_1110001_0000010_1101011;
  end
endmodule
